`define Instset_Wid    63

`define Zero_Word      32'b0

`define F_D_Wid        35
`define Bran_Wid       33
`define D_E_Wid        313
`define E_M_Wid        224+32
`define M_W_Wid        136

`define E_RF_Wid       104
`define M_RF_Wid       104
`define W_RF_Wid       104
`define HILO_Wid       66

`define CP0_Reg_badaddr     5'b01000
`define CP0_Reg_status      5'b01100
`define CP0_Reg_cause       5'b01101 
`define CP0_Reg_epc         5'b01110
`define CP0_Reg_count       5'b01001
`define CP0_Reg_compare     5'b01011

